package alu_pkg;
  `include "transaction.sv"
  `include "generator.sv"
  `include "driver.sv"
  `include "reference_model.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "test.sv"
endpackage
~
