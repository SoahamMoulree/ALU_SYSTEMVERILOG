`define no_of_testcases 500
`define W 8
`define N 4
`define SHIFT_WIDTH  $clog2(`W)
